
module S_P (
	probe,
	source);	

	input	[255:0]	probe;
	output	[255:0]	source;
endmodule
